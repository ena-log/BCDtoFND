`timescale 1ns / 1ps

module FND_SelectDecoder(
    //input, output?? wire type
    input [1:0] i_digitSelect,
    input i_en,                 //enable
    output [3:0] o_digit
    );

    //reg type : memory ???
    reg [3:0] r_digit;
    assign o_digit = r_digit;

    // always @() : ?????? ?????? ???????? ???? ????????? ???????
    // -> always @(i_digitSelect) : ?????? ????????? ???? ??????
    // (i_digitSelect, i_en) == (i_digitSelect or i_en)
    always @(i_digitSelect, i_en) begin
        // if else ???? always ??????????? ??? ??? ??????
        if (i_en) begin
            r_digit = 4'b1111;
        end
        else begin
            case (i_digitSelect)            // c?????? swich ????
                2'h0 : r_digit = 4'b1110;   // c?????? case ????
                2'h1 : r_digit = 4'b1101;
                2'h2 : r_digit = 4'b1011;
                2'h3 : r_digit = 4'b0111;
            endcase
        end
    end

endmodule
